
// Discription: APB Interface
interface apb_interface(input pclk,prst);

endinterface
