`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "ahb_transaction.sv"
`include "ahb_interface.sv"
`include "ahb_driver.sv"
`include "ahb_sequencer.sv"
`include "ahb_monitor.sv"
`include "ahb_coverage.sv"
`include "ahb_responder.sv"
`include "ahb_agent.sv"
`include "ahb_env.sv"
`include "ahb_base_test.sv"
`include "ahb_top.sv"