`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "apb_base_test.sv"
`include "apb_env.sv"
`include "apb_agent.sv"
`include "apb_driver.sv"
`include "apb_sequencer.sv"
`include "apb_monitor.sv"
`include "apb_coverage.sv"
`include "apb_rsponder.sv"
`include "apb_transaction.sv"
`include "apb_top.sv"
