// Discription: AHB Sequencer

typedef uvm_sequencer#(ahb_transaction) ahb_sequencer; 
