interface ahb_interface(input clk,rst);

endinterface
