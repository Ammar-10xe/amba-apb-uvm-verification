
class ahb_transaction extends uvm_sequence_item;
        `uvm_object_utils(ahb_transaction);

        function new(string name = "");
                super.new(name);
        endfunction

        
        
endclass
