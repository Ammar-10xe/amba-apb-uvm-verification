// Discription: APB Sequencer

typedef uvm_sequencer#(apb_transaction) apb_sequencer; 
