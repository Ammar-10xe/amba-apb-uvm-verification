// Discription: axi Sequencer

typedef uvm_sequencer#(axi_transaction) axi_sequencer; 
