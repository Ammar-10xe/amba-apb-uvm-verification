`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "axi_transaction.sv"
`include "axi_interface.sv"
`include "axi_driver.sv"
`include "axi_sequencer.sv"
`include "axi_monitor.sv"
`include "axi_coverage.sv"
`include "axi_responder.sv"
`include "axi_agent.sv"
`include "axi_env.sv"
`include "axi_scoreboard.sv"
`include "axi_base_test.sv"
`include "axi_top.sv"
